LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY tb_transceiverFSMControl IS
END tb_transceiverFSMControl;

ARCHITECTURE behavior OF tb_transceiverFSMControl IS

  -- Component Declaration
  COMPONENT transceiverFSMControl
    PORT(
      TDRE, TSRF, TXD, C8 : IN  STD_LOGIC;
      G_Clock             : IN  STD_LOGIC;
      G_Reset             : IN  STD_LOGIC;
      resetCount          : OUT STD_LOGIC;
      shiftEN             : OUT STD_LOGIC;
      loadEN              : OUT STD_LOGIC;
      TXOut               : OUT STD_LOGIC;
      stateOut            : OUT STD_LOGIC_VECTOR(2 downto 0)
    );
  END COMPONENT;

  -- Constants
  CONSTANT clock_period : TIME := 10 ns;

  -- Input Signals
  SIGNAL TDRE     : STD_LOGIC := '1';
  SIGNAL TSRF     : STD_LOGIC := '0';
  SIGNAL TXD      : STD_LOGIC := '0';
  SIGNAL C8       : STD_LOGIC := '0';
  SIGNAL G_Clock  : STD_LOGIC := '0';
  SIGNAL G_Reset  : STD_LOGIC := '0';

  -- Output Signals
  SIGNAL resetCount : STD_LOGIC;
  SIGNAL shiftEN    : STD_LOGIC;
  SIGNAL loadEN     : STD_LOGIC;
  SIGNAL TXOut      : STD_LOGIC;
  SIGNAL stateOut   : STD_LOGIC_VECTOR(2 downto 0);

  -- Clock control
  SIGNAL stop_clock : BOOLEAN := FALSE;

  -- State constants for readability
  CONSTANT STATE_A : STD_LOGIC_VECTOR(2 downto 0) := "000";  -- Idle
  CONSTANT STATE_B : STD_LOGIC_VECTOR(2 downto 0) := "001";  -- Load
  CONSTANT STATE_C : STD_LOGIC_VECTOR(2 downto 0) := "010";  -- Shift1
  CONSTANT STATE_D : STD_LOGIC_VECTOR(2 downto 0) := "011";  -- Shift2
  CONSTANT STATE_E : STD_LOGIC_VECTOR(2 downto 0) := "100";  -- Done

  -- Helper function to convert state to string
  FUNCTION state_to_string(s : STD_LOGIC_VECTOR(2 downto 0)) RETURN STRING IS
  BEGIN
    CASE s IS
      WHEN "000" => RETURN "sA (Idle)";
      WHEN "001" => RETURN "sB (Load)";
      WHEN "010" => RETURN "sC (Shift1)";
      WHEN "011" => RETURN "sD (Shift2)";
      WHEN "100" => RETURN "sE (Done)";
      WHEN OTHERS => RETURN "UNKNOWN";
    END CASE;
  END FUNCTION;

BEGIN

  -- Instantiate the Unit Under Test (UUT)
  uut: transceiverFSMControl
    PORT MAP(
      TDRE       => TDRE,
      TSRF       => TSRF,
      TXD        => TXD,
      C8         => C8,
      G_Clock    => G_Clock,
      G_Reset    => G_Reset,
      resetCount => resetCount,
      shiftEN    => shiftEN,
      loadEN     => loadEN,
      TXOut      => TXOut,
      stateOut   => stateOut
    );

  -- Clock Generation Process
  clock_process: PROCESS
  BEGIN
    WHILE NOT stop_clock LOOP
      G_Clock <= '0';
      WAIT FOR clock_period/2;
      G_Clock <= '1';
      WAIT FOR clock_period/2;
    END LOOP;
    WAIT;
  END PROCESS;

  -- Stimulus Process
  stim_proc: PROCESS
    VARIABLE test_passed : INTEGER := 0;
    VARIABLE test_failed : INTEGER := 0;
  BEGIN
    REPORT "========================================";
    REPORT "Starting transceiverFSMControl Testbench";
    REPORT "========================================";

    -- Test 1: Asynchronous Reset
    REPORT "Test 1: Asynchronous Reset (G_Reset = '0')";
    G_Reset <= '0';
    TDRE <= '1';
    TSRF <= '0';
    TXD <= '0';
    C8 <= '0';
    WAIT FOR clock_period * 2;
    
    IF stateOut = STATE_A THEN
      REPORT "  PASS: Reset to State A (Idle)";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: Expected State A, got " & state_to_string(stateOut) SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    IF TXOut = '1' THEN
      REPORT "  PASS: TXOut = '1' in State A";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: TXOut should be '1' in State A" SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    -- Release reset
    G_Reset <= '1';
    WAIT FOR clock_period;

    -- Test 2: Stay in State A when TDRE = '1'
    REPORT "Test 2: Stay in State A (TDRE = '1')";
    TDRE <= '1';
    WAIT FOR clock_period * 2;
    WAIT FOR 1 ns;
    
    IF stateOut = STATE_A THEN
      REPORT "  PASS: Remained in State A";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: Should remain in State A" SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    -- Test 3: Transition from State A to State B (TDRE = '0')
    REPORT "Test 3: Transition A -> B (TDRE = '0')";
    TDRE <= '0';
    WAIT FOR clock_period;
    WAIT FOR 1 ns;
    
    IF stateOut = STATE_B THEN
      REPORT "  PASS: Transitioned to State B";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: Expected State B, got " & state_to_string(stateOut) SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    IF loadEN = '1' THEN
      REPORT "  PASS: loadEN = '1' in State B";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: loadEN should be '1' in State B" SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    -- Test 4: Stay in State B when TSRF = '0'
    REPORT "Test 4: Stay in State B (TSRF = '0')";
    TSRF <= '0';
    WAIT FOR clock_period;
    WAIT FOR 1 ns;
    
    IF stateOut = STATE_B THEN
      REPORT "  PASS: Remained in State B";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: Should remain in State B" SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;


    -- Test 5: Transition from State B to State C (TSRF = '1')
    REPORT "Test 5: Transition B -> C (TSRF = '1')";
    TSRF <= '1';
    WAIT FOR clock_period;
    WAIT FOR 1 ns;
    
    IF stateOut = STATE_C THEN
      REPORT "  PASS: Transitioned to State C";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: Expected State C, got " & state_to_string(stateOut) SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    IF shiftEN = '1' THEN
      REPORT "  PASS: shiftEN = '1' in State C";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: shiftEN should be '1' in State C" SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;



        -- Test 6: Stay in State C when TXD = '1'
    REPORT "Test 6: Stay in State C (TXD = '1')";
    TXD <= '1';
    WAIT FOR clock_period;
    WAIT FOR 1 ns;
    
    IF stateOut = STATE_C THEN
      REPORT "  PASS: Remained in State C";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: Should remain in State C" SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    -- Test 7: Transition from State C to State D (TXD = '0')
    REPORT "Test 7: Transition C -> D (TXD = '0')";
    TXD <= '0';
    WAIT FOR clock_period;
    WAIT FOR 1 ns;
    
    IF stateOut = STATE_D THEN
      REPORT "  PASS: Transitioned to State D";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: Expected State D, got " & state_to_string(stateOut) SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    IF shiftEN = '1' THEN
      REPORT "  PASS: shiftEN = '1' in State D";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: shiftEN should be '1' in State D" SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    -- Test 8: Stay in State D when C8 = '0'
    REPORT "Test 8: Stay in State D (C8 = '0')";
    C8 <= '0';
    WAIT FOR clock_period * 2;
    WAIT FOR 1 ns;
    
    IF stateOut = STATE_D THEN
      REPORT "  PASS: Remained in State D";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: Should remain in State D" SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    -- Test 9: Transition from State D to State E (C8 = '1')
    REPORT "Test 9: Transition D -> E (C8 = '1')";
    C8 <= '1';
    WAIT FOR clock_period;
    WAIT FOR 1 ns;
    
    IF stateOut = STATE_E THEN
      REPORT "  PASS: Transitioned to State E";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: Expected State E, got " & state_to_string(stateOut) SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    IF TXOut = '1' THEN
      REPORT "  PASS: TXOut = '1' in State E";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: TXOut should be '1' in State E" SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    -- Test 10: Stay in State E when TDRE = '1'
    REPORT "Test 10: Stay in State E (TDRE = '1')";
    TDRE <= '1';
    WAIT FOR clock_period * 2;
    WAIT FOR 1 ns;
    
    IF stateOut = STATE_E THEN
      REPORT "  PASS: Remained in State E";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: Should remain in State E" SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    -- Test 11: Transition from State E to State A (TDRE = '0')
    REPORT "Test 11: Transition E -> A (TDRE = '0')";
    TDRE <= '0';
    WAIT FOR clock_period;
    WAIT FOR 1 ns;
    
    IF stateOut = STATE_A THEN
      REPORT "  PASS: Transitioned back to State A";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: Expected State A, got " & state_to_string(stateOut) SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    -- Test 12: Full cycle test
    REPORT "Test 12: Complete State Cycle";
    TDRE <= '1';
    TSRF <= '0';
    TXD <= '0';
    C8 <= '0';
    WAIT FOR clock_period;  -- Should stay in A
    
    TDRE <= '0';
    WAIT FOR clock_period;  -- A -> B
    WAIT FOR 1 ns;
    IF stateOut = STATE_B THEN
      test_passed := test_passed + 1;
    ELSE
      test_failed := test_failed + 1;
    END IF;
    
    TSRF <= '1';
    WAIT FOR clock_period;  -- B -> C
    WAIT FOR 1 ns;
    IF stateOut = STATE_C THEN
      test_passed := test_passed + 1;
    ELSE
      test_failed := test_failed + 1;
    END IF;
    
    TXD <= '0';
    WAIT FOR clock_period;  -- C -> D
    WAIT FOR 1 ns;
    IF stateOut = STATE_D THEN
      test_passed := test_passed + 1;
    ELSE
      test_failed := test_failed + 1;
    END IF;
    
    C8 <= '1';
    WAIT FOR clock_period;  -- D -> E
    WAIT FOR 1 ns;
    IF stateOut = STATE_E THEN
      test_passed := test_passed + 1;
    ELSE
      test_failed := test_failed + 1;
    END IF;
    
    TDRE <= '0';
    WAIT FOR clock_period;  -- E -> A
    WAIT FOR 1 ns;
    IF stateOut = STATE_A THEN
      REPORT "  PASS: Complete cycle successful";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: Cycle did not complete correctly" SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    -- Test 13: Reset during active operation
    REPORT "Test 13: Reset During Operation";
    TDRE <= '0';
    WAIT FOR clock_period * 2;  -- Move to State B
    G_Reset <= '0';
    WAIT FOR clock_period;
    WAIT FOR 1 ns;
    
    IF stateOut = STATE_A THEN
      REPORT "  PASS: Reset during operation works";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: Reset failed during operation" SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;
    
    G_Reset <= '1';
    WAIT FOR clock_period;

    -- Test 14: resetCount signal check
    REPORT "Test 14: resetCount Signal";
    TDRE <= '0';
    TSRF <= '0';
    WAIT FOR clock_period;  -- Go to State B
    WAIT FOR 1 ns;
    
    -- resetCount should be asserted in next cycle when in B and w=1
    TSRF <= '1';  -- This makes w=1 in state B
    WAIT FOR clock_period;
    WAIT FOR 1 ns;
    
    IF resetCount = '1' THEN
      REPORT "  PASS: resetCount asserted correctly";
      test_passed := test_passed + 1;
    ELSE
      REPORT "  FAIL: resetCount not asserted" SEVERITY ERROR;
      test_failed := test_failed + 1;
    END IF;

    -- Final Summary
    REPORT "========================================";
    REPORT "Testbench Completed";
    REPORT "========================================";
    
    IF test_failed = 0 THEN
      REPORT "*** ALL TESTS PASSED ***" SEVERITY NOTE;
    ELSE
      REPORT "*** SOME TESTS FAILED ***" SEVERITY ERROR;
    END IF;
    
    REPORT "========================================";
    
    stop_clock <= TRUE;
    WAIT;
  END PROCESS;

END behavior;
